
--defining nand
entity nand_gate is
	Port (a : in std_logic; b: in std_logic; f: in std_logic);
end nand_gate;


	
	